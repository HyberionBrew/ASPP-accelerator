LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

USE work.core_pck.ALL;
USE IEEE.math_real.ALL;

PACKAGE control_pck IS

	CONSTANT DEPTH_PSUM_BUFFER : NATURAL := IFMAP_SIZE * (IFMAP_SIZE/PE_COLUMNS); --33*11
	CONSTANT AWIDTH_PSUM_BUFFER : NATURAL := INTEGER(ceil(log2(real(DEPTH_PSUM_BUFFER))));
	CONSTANT DWIDTH_PSUM_BUFFER : NATURAL := PARALLEL_OFMS * ACC_DATA_WIDTH * PE_COLUMNS;


	CONSTANT AWIDTH_IACTS_BUFFER: NATURAL := INTEGER(ceil(log2(real(FILTER_DEPTH * IFMAP_SIZE * IFMAP_SIZE * 2))));
	CONSTANT DEPTH_IACTS_BUFFER: NATURAL := FILTER_DEPTH * 2 * IFMAP_SIZE * IFMAP_SIZE;
	
	TYPE iacts_buffer_type IS ARRAY(0 TO PE_COLUMNS - 1, 0 TO FILTER_PER_PE - 1) OF unsigned(DATA_WIDTH - 1 DOWNTO 0);
	TYPE array_buffer IS ARRAY(0 TO 36 - 1) OF unsigned(DATA_WIDTH - 1 DOWNTO 0);
	TYPE iacts_mode_type IS (ENABLE_MEM, LOAD_IFMAP, PREPARE_IFMAP, CLEAN);
	TYPE mode_psums_type IS (PREPARE_PSUMS, FETCH_PSUMS, WRITE_BACK, CLEAN, WRITE_OUT_PSUMS);

	TYPE ifmap_address_type IS RECORD
		shared_address : NATURAL;
		shared_address_offset : NATURAL RANGE 0 TO 8;
		address : NATURAL;
	END RECORD;

	TYPE psum_address_type IS RECORD
		x : NATURAL RANGE 0 TO IFMAP_SIZE/PE_COLUMNS - 1;
		y : NATURAL RANGE 0 TO IFMAP_SIZE - 1;
		ofm : NATURAL RANGE 0 TO 3 - 1; --not used->because in parallel TODO! check
	END RECORD;

	TYPE ifmap_position_type IS RECORD
		x : NATURAL RANGE 0 TO IFMAP_SIZE/PE_COLUMNS - 1;
		y : NATURAL RANGE 0 TO IFMAP_SIZE - 1;
		depth_pos : NATURAL RANGE 0 TO FILTER_DEPTH - 1;
	END RECORD;

	TYPE point IS RECORD
		x : NATURAL RANGE 0 TO IFMAP_SIZE/PE_COLUMNS - 1;
		y : NATURAL RANGE 0 TO IFMAP_SIZE - 1;
	END RECORD;

	FUNCTION to_buffer(v : STD_LOGIC_VECTOR(144 * 2 - 1 DOWNTO 0)) RETURN array_buffer;

END PACKAGE;

PACKAGE BODY control_pck IS
	FUNCTION to_buffer(v : STD_LOGIC_VECTOR(144 * 2 - 1 DOWNTO 0)) RETURN array_buffer IS
		VARIABLE buf : array_buffer := (OTHERS => (OTHERS => '0'));
	BEGIN
		FOR I IN 0 TO 36 - 1 LOOP
			buf(I) := unsigned(v(DATA_WIDTH * (I + 1) - 1 DOWNTO DATA_WIDTH * I));
		END LOOP;
		RETURN buf;
	END FUNCTION;

END PACKAGE BODY;
