LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.core_pck.ALL;

PACKAGE pe_pack IS
  CONSTANT COMPARISON_BITVEC_WIDTH : NATURAL := 16;
  CONSTANT DATA_WIDTH_RESULT : NATURAL := 18;
END PACKAGE;