LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE core_pck IS
  CONSTANT FILTER_DEPTH : NATURAL := 10;
  CONSTANT PARALLEL_OFMS : NATURAL := 32;
  CONSTANT MAX_OFMS : NATURAL := 32;
  CONSTANT PE_COLUMNS : NATURAL := 3;
  CONSTANT OFM_REQUANT : NATURAL := 66;
  CONSTANT IFMAP_ZERO_CONSTANT : NATURAL := 24;
  CONSTANT DATA_WIDTH : NATURAL := 8;
  CONSTANT FILTER_PER_PE : NATURAL := 64;
  CONSTANT BUSSIZE : NATURAL := FILTER_PER_PE * DATA_WIDTH + FILTER_PER_PE; -- data +bitvec + ifmap zero offset + Ifmap_zero
  CONSTANT MAX_RATE : NATURAL := 1;
  CONSTANT ACC_DATA_WIDTH : NATURAL := 24;
  CONSTANT EXEC_COUNTER_WIDTH : NATURAL := 32;
  
  CONSTANT IFMAP_SIZE : NATURAL := 33;
  CONSTANT DILATION_RATE : NATURAL := 6;

END PACKAGE;